//----------------------------------------------------------------------------
//-- Declare machine cycle and instruction cycle parameters
//----------------------------------------------------------------------------

// RV32I Base Integer Instructions

localparam [6:0] lw 
